acl:attr
acl:relat
advmod:emph
aux:neg
flat:foreign
flat:name
nmod:attr
nmod:poss
nmod:relat
parataxis:speech
