acl:att
acl:av
acl:cleft
acl:efter
acl:från
acl:för
acl:hos
acl:huruvida
acl:i
acl:innan
acl:liksom
acl:med
acl:mot
acl:när
acl:om
acl:på
acl:relcl
acl:som
acl:såsom
acl:till
acl:utan
acl:vid
acl:än
acl:över
advcl:allt_efter_som
advcl:allt_eftersom
advcl:alltefter_som
advcl:allteftersom
advcl:antingen
advcl:att
advcl:av
advcl:beroende_på
advcl:bortsett_från
advcl:dess
advcl:därför_att
advcl:då
advcl:då_och_då
advcl:efter
advcl:efter_att
advcl:efter_det_att
advcl:efter_hand_som
advcl:eftersom
advcl:ehuruväl
advcl:emedan
advcl:fast
advcl:fastän
advcl:från
advcl:från_det
advcl:för
advcl:för_att
advcl:förrän
advcl:förutsatt_att
advcl:genom
advcl:hos
advcl:i
advcl:i_de_fall
advcl:i_samband_med
advcl:i_stället_för
advcl:if
advcl:ifråga_om
advcl:innan
advcl:liksom
advcl:låt_vara
advcl:med
advcl:medan
advcl:när
advcl:nära
advcl:oavsett
advcl:oberoende_av
advcl:om
advcl:på
advcl:på_det
advcl:samtidigt_med_att
advcl:samtidigt_som
advcl:sedan
advcl:som
advcl:så
advcl:så_att
advcl:så_fort
advcl:så_länge
advcl:så_långt
advcl:så_snart
advcl:såsom
advcl:såvida
advcl:till
advcl:tills
advcl:trots_att
advcl:under_det_att
advcl:under_förutsättning_att
advcl:utan
advcl:utöver
advcl:vare_sig
advcl:än
advcl:även_om
advcl:över
aux:pass
compound:prt
conj:and
conj:el
conj:eller
conj:fast
conj:för
conj:men
conj:och
conj:plus
conj:resp
conj:respektive
conj:samt
conj:som
conj:sym
conj:så
conj:såväl_som
conj:ty
conj:utan
csubj:pass
flat:name
nmod:a
nmod:angående
nmod:av
nmod:bak
nmod:bakom
nmod:beträffande
nmod:bland
nmod:bredvid
nmod:de
nmod:efter
nmod:emellan
nmod:enligt
nmod:f
nmod:for
nmod:fr_o_m
nmod:framför
nmod:från
nmod:för
nmod:för_sedan
nmod:före
nmod:genom
nmod:gentemot
nmod:hos
nmod:i
nmod:i_form_av
nmod:i_fråga_om
nmod:i_förening_med
nmod:i_förhållande_till
nmod:i_linje_med
nmod:i_proportion_till
nmod:i_samarbete_med
nmod:i_samband_med
nmod:in
nmod:inför
nmod:inklusive
nmod:inom
nmod:intill
nmod:jämfört_med
nmod:jämte
nmod:kontra
nmod:kring
nmod:längs
nmod:med
nmod:med_avseende_på
nmod:med_hjälp_av
nmod:med_hänsyn_till
nmod:med_sikte_på
nmod:mellan
nmod:mot
nmod:när_det_gällde
nmod:när_det_gäller
nmod:nära
nmod:oavsett
nmod:of
nmod:om
nmod:omkring
nmod:ovanför
nmod:ovanpå
nmod:per
nmod:plus
nmod:poss
nmod:på
nmod:på_grund
nmod:på_grund_av
nmod:runt
nmod:rörande
nmod:sedan
nmod:sym
nmod:t_o_m
nmod:till
nmod:till_förmån_för
nmod:under
nmod:ur
nmod:utan
nmod:utanför
nmod:utom
nmod:utöver
nmod:vad_gäller
nmod:via
nmod:vid
nmod:vid_sidan_om
nmod:à
nmod:åt
nmod:över
nsubj:pass
obl:agent
obl:allt_efter
obl:alltefter
obl:av
obl:bakom
obl:beroende_på
obl:beträffande
obl:bland
obl:bortsett_från
obl:efter
obl:emellan
obl:emot
obl:enl
obl:enligt
obl:exkl
obl:fr_o_m
obl:framemot
obl:framför
obl:from
obl:från
obl:från_och_med
obl:frånsett
obl:för
obl:för_sedan
obl:för_sen
obl:för_skull
obl:förbi
obl:före
obl:förrän
obl:förutan
obl:förutom
obl:genom
obl:gentemot
obl:hos
obl:i
obl:i_anslutning_till
obl:i_enlighet_med
obl:i_form_av
obl:i_fråga_om
obl:i_förbindelse_med
obl:i_förhållande_till
obl:i_jämförelse_med
obl:i_motsats_till
obl:i_mån_av
obl:i_närheten_av
obl:i_och_med
obl:i_proportion_till
obl:i_riktning_mot
obl:i_samband_med
obl:i_skydd_av
obl:i_stället_för
obl:i_takt_med
obl:ifråga_om
obl:ifrån
obl:igenom
obl:inför
obl:innanför
obl:inom
obl:inom_ramen_för
obl:inpå
obl:intill
obl:istället_för
obl:jämfört_med
obl:kring
obl:liksom
obl:längs
obl:lågstadiet
obl:med
obl:med_avseende_på
obl:med_hjälp_av
obl:med_hänsyn_till
obl:med_hänvisning_till
obl:med_tanke_på
obl:med_undantag_för
obl:med_utgångspunkt_av
obl:med_utgångspunkt_i
obl:mellan
obl:mot
obl:nedanför
obl:nedom
obl:när_det_gällde
obl:när_det_gäller
obl:när_det_gällt
obl:nära
obl:närmare
obl:oavsett
obl:oberoende_av
obl:om
obl:omkring
obl:ovanför
obl:ovanpå
obl:over
obl:per
obl:på
obl:på_basis_av
obl:på_grund_av
obl:på_grundval_av
obl:på_tal_om
obl:på_tredje
obl:runt
obl:runtomkring
obl:sedan
obl:senast
obl:som
obl:sym
obl:t_o_m
obl:tack_vare
obl:tidigast
obl:till
obl:till_följd_av
obl:till_höger_om
obl:till_skillnad_från
obl:till_skillnad_mot
obl:till_vänster_om
obl:tom
obl:trots
obl:tvärsigenom
obl:tvärtemot
obl:under
obl:under_loppet_av
obl:ur
obl:utan
obl:utan_avseende_på
obl:utan_hänsyn_till
obl:utan_tanke_på
obl:utanför
obl:utifrån
obl:utom
obl:utåt
obl:utöver
obl:vad_beträffar
obl:vad_det_gäller
obl:vad_gäller
obl:via
obl:vid
obl:vid_sidan_av
obl:vid_sidan_om
obl:värld
obl:än
obl:å
obl:åt
obl:över
