VerbForm=Stem
