nmod:poss
acl:relcl
compound:prt
nmod:agent
