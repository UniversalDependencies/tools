advcl:om
nmod:av
nmod:i
nmod:på
obl:agent:av
obl:av
obl:i
obl:på
