acl:relcl
compound:prt
nmod:agent
nmod:poss
