acl:relcl
compound:prt
nmod:poss
obl:agent
