[B|b]l a
[D|d] v s
[E|e] d
[F|f] n
[F|f]r o m
[M|m] fl
[M|m] m
[O|o] s v
[S|s] k
[T|t] ex
[T|t] o m
[T|t] v
