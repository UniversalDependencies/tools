advcl:att
advcl:då
advcl:efter_det_att
advcl:eftersom
advcl:för_att
advcl:förutsatt_att
advcl:innan
advcl:liksom
advcl:medan
advcl:när
advcl:oavsett
advcl:om
advcl:på
advcl:utan
advcl:sedan
advcl:som
advcl:så_att
advcl:såsom
advcl:utan
advcl:även_om
nmod:av
nmod:i
nmod:plus
nmod:på
obl:agent:av
obl:av
obl:för
obl:i
obl:med
obl:på
obl:till
