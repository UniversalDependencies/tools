acl:cleft
acl:relcl
aux:pass
compound:prt
csubj:pass
flat:name
nmod:poss
nsubj:pass
obl:agent
