[Bb]l a
[Dd] v s
[Ee] d
[Ff] n
[Ff]r o m
[Mm] fl
[Mm] m
[Oo] s v
[Ss] k
[Tt] ex
[Tt] o m
[Tt] v
